`include "ingle_Cycle_Top"

module top();











endmodule